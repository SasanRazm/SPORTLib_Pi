.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=120OHM, RN=14OHM, ICRIT=0.6MA)
.MODEL PIJJ JJ(RTYPE=1, VG=2.8MV, CAP=0.04PF, R0=20OHM, RN=8OHM, ICRIT=1MA, PHI=PI)

.subckt JTL 1 9
L1 1 2 0.1p

B1 2 12 PIJJ area=0.03
Lpi 12 0 0.3pH

LP2 2 3 0.15pH
B2 3 4 JJMIT area=0.07
LP3 4 5 0.15pH
B3 5 6 JJMIT area=0.07
LP4 6 7 0.15pH
B4 7 8 JJMIT area=0.07
LP5 8 9 0.15pH

IB1 0 2 pwl(0 0 10ps 15uA)
.ends

.SUBCKT DCSFQ 1 13
L1 2 3 0.1p
RINON 1 2 50OHM
LGND 2 0  1pH

BIN 3 4 JJMIT area=0.08
LPIN 4 5 0.1pH

B1 5 6 PIJJ area=0.03
Lpi 6 0 0.3pH

LP2 5 7 0.1pH
B2 7 8 JJMIT area=0.07
LP3 8 9 0.1pH
B3 9 10 JJMIT area=0.07
LP4 10 11 0.1pH
B4 11 12 JJMIT area=0.07
LP5 12 13 0.1pH

IB1 0 5 pwl(0 0 10ps 10uA)
.ends

.SUBCKT DFF 1 21 16

LP1 1 2 0.2p
B1 2 0 PIJJ AREA=0.03

LP2 2 3 0.1pH
B2 3 4 JJMIT area=0.075
LP3 4 5 0.1pH
B3 5 6 PIJJ area=0.03
LP4 6 9 0.1pH


B5 9 0 PIJJ AREA=0.03

LPCLK 21 22 0.2p
B6 22 9 JJMIT AREA=0.05

B7 9 10 JJMIT area=0.09
LP6 10 11 0.1pH
B8 11 12 JJMIT area=0.09
LP7 12 13 0.1pH
B9 13 14 JJMIT area=0.09
LP8 14 15 0.1pH

LPOUT 15 16 0.2p

IB1 0 2 pwl(0 0 10ps 10uA)
IB2 0 9 pwl(0 0 10ps 20uA)
.ENDS DFF

X11 DCSFQ 22 1
X1 JTL 1 2
X2 JTL 2 3
X3 JTL 3 4
X4 JTL 4 5

X44 DCSFQ 44 6
X5 JTL 6 7
X6 JTL 7 8
X7 JTL 8 9
X8 JTL 9 10

X9 DFF 5 10 11
X10 JTL 11 12
X12 JTL 12 13

V1 22 0 PULSE(0.0mv  30mv   230ps   3.0ps   3.0ps   5.0ps   40.0ps)
V2 44 0 PULSE(0.0mv  30mv   20ps   3.0ps   3.0ps   5.0ps   20.0ps)

Lload 13 17 5pH
RNONload 17 0 50ohm

.TRAN 0.1PS 600PS 500PS 0.1PS
.FILE OUT.CSV
.PRINT NODEV 5 0
.PRINT NODEV 10 0
.PRINT NODEV 11 0
