.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=120OHM, RN=14OHM, ICRIT=0.6MA)
.MODEL PIJJ JJ(RTYPE=1, VG=2.8MV, CAP=0.04PF, R0=20OHM, RN=8OHM, ICRIT=1MA, PHI=PI)

.subckt JTL 1 9
L1 1 2 0.1p

B1 2 12 PIJJ area=0.03
Lpi 12 0 0.3pH

LP2 2 3 0.15pH
B2 3 4 JJMIT area=0.07
LP3 4 5 0.15pH
B3 5 6 JJMIT area=0.07
LP4 6 7 0.15pH
B4 7 8 JJMIT area=0.07
LP5 8 9 0.15pH

IB1 0 2 pwl(0 0 10ps 15uA)
.ends

XIN 23 1 JTL
X1 1 2 JTL
X2 2 3 JTL
X3 3 4 JTL
X4 4 5 JTL
X5 5 6 JTL
X6 6 7 JTL
X7 7 8 JTL
X8 8 9 JTL
X9 9 10 JTL
X10 10 11 JTL
X11 11 12 JTL
X12 12 13 JTL
X13 13 14 JTL
X14 14 15 JTL
X15 15 16 JTL
Lload 16 17 5pH
RNONload 17 0 50ohm

V1 23  22 PULSE(0.0mv  0.6mv   50ps   2.0ps   2.0ps   1.0ps   10.0ps)
RNONIN 0 22 10ohm

.tran 0.025p 1000p 950p 0.025p
.FILE OUT.CSV
.print nodev 6 0
*.print nodev 11 0
.print nodev 16 0
