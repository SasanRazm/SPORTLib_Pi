.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=120OHM, RN=14OHM, ICRIT=0.6MA)
.MODEL PIJJ JJ(RTYPE=1, VG=2.8MV, CAP=0.04PF, R0=20OHM, RN=8OHM, ICRIT=1MA, PHI=PI)

.subckt JTL 1 9
L1 1 2 0.1p

B1 2 12 PIJJ area=0.03
Lpi 12 0 0.3pH

LP2 2 3 0.15pH
B2 3 4 JJMIT area=0.07
LP3 4 5 0.15pH
B3 5 6 JJMIT area=0.07
LP4 6 7 0.15pH
B4 7 8 JJMIT area=0.07
LP5 8 9 0.15pH

IB1 0 2 pwl(0 0 10ps 15uA)
.ends

.SUBCKT DCSFQ 1 13
L1 2 3 0.1p
RINON 1 2 50OHM
LGND 2 0  1pH

BIN 3 4 JJMIT area=0.08
LPIN 4 5 0.1pH

B1 5 6 PIJJ area=0.03
Lpi 6 0 0.3pH

LP2 5 7 0.1pH
B2 7 8 JJMIT area=0.07
LP3 8 9 0.1pH
B3 9 10 JJMIT area=0.07
LP4 10 11 0.1pH
B4 11 12 JJMIT area=0.07
LP5 12 13 0.1pH

IB1 0 5 pwl(0 0 10ps 10uA)
.ends

.subckt JTLs 1 9
L1 1 2 0.1p
B1 2 12 PIJJ area=0.027
Lpi 12 0 0.3pH
LP2 2 3 0.1pH
B2 3 4 JJMIT area=0.065
LP3 4 5 0.1pH
B3 5 6 JJMIT area=0.065
LP4 6 7 0.1pH
B4 7 8 JJMIT area=0.065
LP5 8 9 0.1pH
IB1 0 2 pwl(0 0 10ps 15uA)
.ends

.subckt SPL 1 20 21
L1 1 2 0.1p
B1 2 22 PIJJ area=0.03
Lpi 22 0 0.3pH
LP2 2 3 0.1pH
B2 3 8 JJMIT area=0.042
X1 JTLs 8 20
LP5 2 9 0.1pH
B5 9 14 JJMIT area=0.042
X2 JTLs 14 21
IB1 0 2 pwl(0 0 10ps 25uA)
.ends


X0 DCSFQ 99 1
X1 JTL 1 2
X2 JTL 2 3
X3 SPL 3 5 6
X4 JTL 5 7
X5 JTL 6 8


Lload1 7 17 5pH
RNONload 17 0 300ohm

Lload2 8 18 5pH
RNONload2 18 0 300ohm

V1 99 0 PULSE(0.0mv  30mv   20ps   3.0ps   3.0ps   10.0ps   40.0ps)

.TRAN 0.01PS 600PS 500PS 0.01PS
.FILE OUT.CSV
.PRINT NODEV 99 0
.PRINT NODEV 7 0
.PRINT NODEV 8 0
