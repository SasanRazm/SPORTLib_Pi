.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=120OHM, RN=14OHM, ICRIT=0.6MA)
.MODEL PIJJ JJ(RTYPE=1, VG=2.8MV, CAP=0.04PF, R0=20OHM, RN=8OHM, ICRIT=1MA, PHI=PI)

.subckt JTL 1 9
L1 1 2 0.1p

B1 2 12 PIJJ area=0.03
Lpi 12 0 0.3pH

LP2 2 3 0.15pH
B2 3 4 JJMIT area=0.07
LP3 4 5 0.15pH
B3 5 6 JJMIT area=0.07
LP4 6 7 0.15pH
B4 7 8 JJMIT area=0.07
LP5 8 9 0.15pH

IB1 0 2 pwl(0 0 10ps 15uA)
.ends

.SUBCKT DCSFQ 1 13
L1 2 3 0.1p
RINON 1 2 50OHM
LGND 2 0  1pH

BIN 3 4 JJMIT area=0.08
LPIN 4 5 0.1pH

B1 5 6 PIJJ area=0.03
Lpi 6 0 0.3pH

LP2 5 7 0.1pH
B2 7 8 JJMIT area=0.07
LP3 8 9 0.1pH
B3 9 10 JJMIT area=0.07
LP4 10 11 0.1pH
B4 11 12 JJMIT area=0.07
LP5 12 13 0.1pH

IB1 0 5 pwl(0 0 10ps 10uA)
.ends

.SUBCKT MERGER 1 9 22

LIN1 1 2 0.1p
B1 2 121 PIJJ AREA=0.033
Lp1 121 0 0.3pH

Lp2 2 3 0.1pH
B2 3 4 JJMIT AREA=0.11
Lp3 4 5 0.1pH
B3 5 6 JJMIT AREA=0.11
Lp4 6 7 0.1pH
B4 7 8 PIJJ AREA=0.025

LIN2 9 10 0.2p
B5 10 101 PIJJ AREA=0.033
Lp5 101 0 0.3pH

Lp6 10 11 0.1pH
B6 11 12 JJMIT AREA=0.11
Lp7 12 13 0.1pH
B7 13 14 JJMIT AREA=0.11
Lp8 14 15 0.1pH
B8 15 8 PIJJ AREA=0.025

LP9 8 16 0.1pH

B10 16 161 PIJJ AREA=0.025
LP10 161 0 0.1pH

Lp11 16 17 0.1pH
B12 17 18 JJMIT AREA=0.08
Lp12 18 19 0.1pH
B13 19 20 JJMIT AREA=0.08
Lp13 20 21 0.1pH
B14 21 22 JJMIT AREA=0.08
 
IB1 0 2 pwl(0 0 10ps 15uA)
IB2 0 10 pwl(0 0 10ps 15uA)
IB3 0 16 pwl(0 0 10ps 27uA)
.ENDS

RNONload 17 0 300ohm
LLoad 15 17 5pH

X11 DCSFQ 11 1
X1 JTL 1 2
X2 JTL 2 3
X44 DCSFQ 44 4
X3 JTL 4 5
X4 JTL 5 6
X7 MERGER 3 6 13
X8 JTL 13 14
X9 JTL 14 115
X10 JTL 115 15
V11 111 0  PULSE(0.0mv  30mv   100ps   3.0ps   3.0ps   20.0ps   120.0ps)
V1 11 111 PULSE(0.0mv  30mv   140ps   3.0ps   3.0ps   20.0ps   120.0ps)
V2 44 0 PULSE(0.0mv  30mv   20ps   3.0ps   3.0ps   20.0ps   80.0ps)

.TRAN 0.1PS 440PS 40PS 0.1PS
.FILE OUT.CSV
.PRINT NODEV 3 0
.PRINT NODEV 6 0
.PRINT NODEV 13 0
